* D:\circuit project\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Tue Jan 29 19:33:16 2019



** Analysis setup **
.tran 0 1000
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
